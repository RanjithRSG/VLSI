class i2c_transaction;
  
  logic scl_pad_i;
  logic scl_pad_o;
  logic scl_padoen_o;
  logic sda_pad_i;
  logic sda_pad_o;
  logic sda_padeon_o;
  logic interrupt_o;
  
endclass
