class transaction;
  
  bit clk;
  rand bit reset;
  bit up_down;
  bit [7:0]count;
  
endclass
