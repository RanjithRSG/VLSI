interface operation;
  
  logic clk;
  logic reset;
  logic up_down;
  logic [7:0]count;
  
endinterface
