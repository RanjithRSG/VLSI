class alu_transaction;
  	
    rand bit [7:0] a, b;
    rand bit [1:0] op;
    bit [7:0] expected_result;

//     function new();
//         super.new();
//     endfunction

//     function void print();
//         $display("ALU Transaction: a=%0h, b=%0h, op=%0h, expected=%0h", a, b, op, expected_result);
//     endfunction
  
endclass
