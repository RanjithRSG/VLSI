class transaction;
  
  rand bit D;
  bit clk;
  rand bit reset;
  bit Q;
  
endclass
