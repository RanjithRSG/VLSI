// Code your design here
module encoder4to2(output X,Y ,input A,B,C,D );
  or(X,A,B);
  or a1(Y,A,C);
endmodule
