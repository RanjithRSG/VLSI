interface operation;
  
  logic D; 
  logic clk;
  logic reset;
  logic Q;
  
endinterface
