class transaction;
  
  rand bit a;
  rand bit b;
  reg sum;
  reg carry;

endclass
