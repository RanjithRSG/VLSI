class transaction;
  
  bit clk;
  rand bit reset;
  reg [7:0] count;
  
endclass
