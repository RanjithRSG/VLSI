class alu_transaction;
  	
    rand bit [7:0] a, b;
    rand bit [1:0] op;
    bit [7:0] expected_result;
  
endclass
