interface operation;
  
  logic clk;
  logic reset;
  logic [7:0] count;
  
endinterface
