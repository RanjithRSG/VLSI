interface operation;
  
  logic clk;
  logic reset;
  logic [8:0]data;
  logic [8:0]addr;
  logic write;
  logic read;
  logic [8:0]dataout;
  
endinterface
